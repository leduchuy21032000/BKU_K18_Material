library verilog;
use verilog.vl_types.all;
entity digitalClock_vlg_vec_tst is
end digitalClock_vlg_vec_tst;
